-- IF Stage test bench
library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity IF_Stage_tb is 
end IF_Stage_tb;

architecture IF_stage_arc of IF_Stage_tb is
  component IF_stage is 
  port
  (
    clk: in std_logic:='0';
    en1,en2: in std_logic :='1';
    PCSrc_D: in std_logic :='0';
    PCBra_D: in std_logic_vector(31 downto 0) :=(others =>'0');
    
    inst_out, PCplus4: out std_logic_vector(31 downto 0):=(others =>'0')
    );
  end component;
  
signal clk: std_logic := '0';
signal PCSrc_D: std_logic := '1';
signal en1,en2: std_logic:='1';
signal PCBra_D: std_logic_vector(31 downto 0) := (others=>'0');
signal inst_out,PCplus4: std_logic_vector(31 downto 0):=(others=>'0');

constant clk_period: time:= 100ns;  

begin
uut: IF_Stage
port map(clk=>clk, en1=>en1, en2=>en2, PCSrc_D=>PCSrc_D, 
         PCBra_D=>PCBra_D, inst_out=>inst_out, PCplus4=>PCplus4);
         
 -- clock gen
 clk_process: process

 begin
      clk<='0';
      wait for clk_period/2;
      clk<='1';
      wait for clk_period/2;
    end process;    
 
  stim_proc: process
    begin
      wait for clk_period;
      wait for clk_period;
      PCSrc_D<='0';
    end process;    
  end;
  
      
