-- sign extension block
library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SignExt is 
  port(
    Sin: in std_logic_vector(15 downto 0) ;
    Sout: out std_logic_vector(31 downto 0)
  );
  
end SignExt;

architecture SignExt_a of SignExt is 
begin
  Sout <= X"FFFF" & Sin when Sin(15) ='1' else
  X"0000" & Sin;
end SignExt_a;


